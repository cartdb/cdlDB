







    



    














     














     































  





  











  







































































***************    ************************************************************************************************************************













    





  *****************



















****    ************    ****







    

****

  






















************      ********** 










 


 






    

   ****************************************************************************************************************************************************************************************    ****





 **** ********************************************* *********************************************************************************************************************  *******************  ****************  ****************************  ************









































    








































  





  



****    ********


  


  


       

   

   

   

       



    





  





  





  





  



  



  





  







***************************************************************************************************************************************************************************************************************************************************

  



    





 







     

 


 







     

 


 







    

 


 







 



 


 


 

**************************************************************************************************************************************************************                        






























*****************************************************************************************************************************************************************************************



																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				       																																																																																																																																																																																																																									            					                                																																																																																																																																																																																																																																																																																							                                																																					        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			   																																																																																																																																																			                       										         																																				 																																																																																																																																												 																																																														    																																																																																																																																																																																																																																																																			                        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			     																																																																																																																																																																																																											  																																																																																																																																																																											 																																																																																																																																																																																																																																																										                                                                       																																																																																																																																																											       																																																																																																																																																																																																																																																																																																						   																																																																																																																																													   										   																																																																																																																																																																																																																																																																																																																																																																     																											    																																																																																																																																																	 																																																																																																																																																																																																																																																																																																																						 																																																																																																																																																																																																																																  															  																																																															     																																																																																																																												      																																																																																																																																																																																																											                                                         				 													   									                                                                                                     																																																												                                                                                                                                                                    ..........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                  ..............................................................................................................................................................................................................................................................................................................................    ..............    ...................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   