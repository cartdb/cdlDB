																																																																																																																																																																																																																																	                																																																											  									               					            			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      																																						                                                                     					   																																																											                  													                                                                    																																																																																																																																																																																																										**************  ********																																																									       																	    																					****************																																																																																																																																												    														   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																                                  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				          							 																																																																																 																																																																																																																																																									 																																																																																																																																																																																																																																																																																													           									    																																							                                                                                 																																																																																																												    																																																																																																																																																																																																																																																																																																																								 				 																																	 																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																											       																																																																																																																																																																																																																																																																																																														      																																																																																																																																																																																																																								                  																																																																													


																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																									 																																																																																																				  																																																																																																																												     																																																																																		
     																																																																																																																																																																																																																																																																																																																																																																									                   																																  																			      																																																										    																																																										   																		                                                   ................                ................                                                             ................                               ......                              ..........................................                                                                      ......                                                                                                                                          ....................................................................................................................................................................                        .........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................  ....................................................................................................................................................................................................   ... .........   .........................    .................................................................................................                        .......  ................................................................................................  ............................................................................................................................... ............................  ....  ................................................                  .....................................................................................................................        .......................................................................................................................................                                                        .................................................................................................................................                                                         ...................                             .....................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  