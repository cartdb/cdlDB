																																																																																																																																																																																																																																	                																																																											  									               					            			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      																																						                                                                     					   																																																				                         													                                                                    																																																																																																																																																																																																										**************  ********																																																									       																	    																					****************																																																																																																																																												    														   																																																																																													                     																																																																																																																																																																																																											                                            																																																																																																																																																																																							                                  																																																																																																																																																																																																																																											           																																							      																																																		       																																																																																															    																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																						          							 																																																																																 																																																																																																																																																									 																																																																																																																																																																																																																																																																																													           									    																																							                                                                                 																																																																																																												    																																																																																																																																																																																																																																																																																																																								 				 																																	 																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			       																																																																																																																																																																																																																																																																	       																																																		                																																																																																																															             																																				      								                                																														      																																																																																																												            																																																																																																                  																																																																													


										                    																																																											                                   																																																																																																	                 																	    																																																																																									     																																																																																																																																															    																																																      																																																																																																																		                                																																																																										   																							  																																																																																																																												     																																																																																		
     																																																																																																																																																																																																																																																																																																																																																																									                   																																  																			      																																																										    																																																					        																		                                                   ................                ................                                                                                                                              ................                                                                                                 ......                                                         ...............                                                                      ......                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ....................................................................................................................................................................                            .....................................................................................................................................................................................................................................................................................................................................................................................................................................................................                ....  .................................................................................................................................................                                      .............   ... ......         ... ........              ......................................                                                                                   .......  ................................................................                                               ...............................................................................................................................    ..............  ..              ..  .....................             ..............                  ............                                                        ..........                   .....................        ......................................................................                   ..............................................                                                                                                                                      ...................................................                                                                                                                                                                                                                                          ...................                             .................................             .......................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  