																																															     																																																																														

















																																																																																																			   																														                    																																					                                        																																																																																																																																																																				     																																																																																																																																									            																																																																													   				   																																																											                                																																																																						

        

        																																												                                                                                                                    																																																																		*******************************************************************************************************************       																																																																																																																																																











																																																													     																																																																																																																																																																																	   
        																																																																																																								  																										



                     



                     																																						           						 																																																																																																		   																																								     																																																																				



 

  

  

  

 
     
     
     
     																																																																																																																																																													   																																																																																																																																				







 

  

  

  

  

  

  

  

  

  

  

  

  








 








 








 

 																																																																																																																																										      															      																																						        				        			 																																																																																													                                              	                                                                                                                                           							                                                                                                                                                                                                                                                                                																                                                                                                                                                                                                                     																																																																																																																														    


















         																																																																					                                                                                                                                                                                                                                                                                                                                                                                                                                                                               																																											
    
    
    
                                                                                                                                                                                                                                                                                                         																																																																																																																																																																																																																																							                                                                                																						     																																																																																																																																																			          






































            
    
        ****                					 	



																																																																	            																																																																																								                                                      																																																																																																																																																																																																																								




											































































































































  																																																																																																																																																											


																																																																																																																																																																																																															








																								




																																																																																																 




 




																																																																															*********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************																																																																			


																															





             


             **********************************                                                                                                                                      *****************                                        ***************************************************************************************************************************************************************                                                                                                               *************************************                                                                                                                                                                   *************************************************                                                                        ********************************                                                                                                                                                    ***************** **********************                                                                **************************                                                                                       ................                                      ............      ........................      ..................      ........................      ......       .........................................................................................................                                   ....................................................................................              ...................................................................................................................................................       ..............                                                                      ..........................................      ..................................................                                                                                                                                                                                                            .....................................                                                                                                    ....                      ........................                       ....................                         ............                                                 ..................................................................................  ...............................................                                                                               ....................................................................                                                                          ....................................................................    .........................                               ............................................................................................................................................................................ .............................................................................................................................................................................................................. ..............................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       