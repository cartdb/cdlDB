																																																																																																																																																																																																																																	                																																																											  									               					            			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      																																						                                                                     					   																																																											                  													                                                                    																																																																																																																																																																																																										**************  ********																																																									       																	    																					****************																																																																																																																																												    														   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																                                  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				          							 																																																																																 																																																																																																																																																																																																																																																																																																																																																																																																																																																							           									    																																							                                                                                 																																																																																																												    																																																																																																																																																																																																																																																																																																																								 				 																																	 																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																											       																																																																																																																																																																																																																																																																																																														      																																																																																																																																																																																																																																		  																																																																																			


																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																									 																																																																																																				  																																																																																																																												     																																																																																		
     																																																																																																																																																																																																																																																																																																																																																																									                   																																  																			      																																																										    																																																										   																		                                                   ................                ................                                          ................                               ......                              ..........................................                                                                      ......                                                                                                                                      ....................................................................................................................................................................                      .........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................  .......................................................................................................................................................................................................... .........   .............................................................................................................................................................  ................................................................................................  ............................................................................................................................... ............................  ....  .......................................................................................................................................................................................        .......................................................................................................................................                                                        .................................................................................................................................                                                         ...................                             .....................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  