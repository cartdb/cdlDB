                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       &&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&                            																								    																																																																																																																				                                            																																																																																								

																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																		 													        																																																																																																																																																																																	  			   


    





    
    






																																																																																																																																																																																																																																																																																																																																																																																																																																																						    																																	                        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																														    																							  																																																												           								                                   																													   																															                             																		       																																  															 																																																	        																																																				                                                                     																																																																                                    																																																									         																												  																																	  																																															                                                      																																																																																				


   																																																********																																																																																																																																																																			  																																																																																																																											       																					  																																			          																														  															                                                                																																																																																																																																																																							    																								                                                              																																																																																																																																																											                																																																																	         																																																																																		                                                                                                                                                                                                                                                                                                                                                                                                                 																																																																		       						                          																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																														  																																																																																																																																																																																																																																																																		                      																																																																																																																																																																																																  																																																																																																																																																																																																					          													                                                                                   																																																																																																******  																																																	  																																																																			                        																		   																																																																														                                                                                       																																																																																																																																																																																																																																																																																																																																																																															  																																		******    ****      **    																																																																																																																																																																																		  																										********************  **    																																																																																			        		             																	                             																				  																																														               			                                                                                              																			  																														    																																																								  																																			                                                                                    																					                         																																																																																							  																																					                     									         																																																																																																		                                                                                ..  ......                                                                                                                                                                                                                                                                                                                                                                                                                                             ........                                                                                                                                                                                                                                                                                                                                                                                                                                                                ..  ..    ..............          ..                                                                                                                     .........                        ......................................................................................................................................................................................                                                                ..............................................                                                                                                                                                 ............................................................................................................................................................                                                                                                                                                                                                                            ............................................................................................................................................................................................................................. ............................................... .........................         ..........................................................................................................................                                                                        .......................                                      ........................................                                                                                ...........................  .........................                         ...........                          .........                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ........          ....................................                                                                                                    ......................................................................                                                            ............................................................................................................................................................................                                                                                                                          ............................................                                  .............................................................................................. . ....... . ....... . ....... . ....... . ....... . ....... . ...... ...... . ...... . ...... . ... . ...... ..... ...... . ...... . .....                                                                                                                                                                                                                                    ....................                                                                                                            ....................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       