                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       &&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&                            																																																																																																																																																                                            																																																																																								

																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																	 													        																																																																																																																																																																																	  			   


    





    
    






																																																																																																																																																																																																																																																																																																																																																																																																																																																						    																																	                        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																														    																							  																																																												           								                                   																																																																							              																									       																																  															 																																																																																																												                                                                     																																																																                                    																																																									         																												  																																	  																																															                                                      																																																																																				


   																																																********																																																																																																																																																																			  																																																																																																																											       																					  																																																																											  															                                                                																																																																																																																																																																							    																								         					        																		         																																																																																																																																																																								                																																																																	         																																																																																		                                                                                                                                                                                                                                                                                                                                                                                                                 																																																																		       																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																														  																																																																																																																																																																																																																																																																		                      																																																																																																																																																																																																  																																																																																																																																																																																																					          													                                                                                   																																																																																																******  																																																	  																																																																			                        																		   																																																																														                                                                                       																																																																																																																																																																																																																																																																																																																																																																															  																																		******    ****      **    																																																																																																																																																																																		  																										********************  **    																																																																																			        		             																	                             																																																																				               			                                                                                              																			  																														    																																																								  																																			                                                                                    																					                         																																																																																																																														                     									         																																																																																																		                                                                                ..  ......                                                                                                                                                                                                                                                                                                                                                                                                                                             ........                                                                                                                                                                                                                                                                                                                                                                                                                                                                ..  ..    ..............          ..                                                                                                                     .........                        ......................................................................................................................................................................................                                                                ..............................................                                                                                                                                                 ............................................................................................................................................................                                                                                                                                                                                                                            ............................................................................................................................................................................................................................. ............................................... .........................         ..........................................................................................................................                                                                        .................................................            ........................................                                                                                ...........................  .........................                         ...........                          .........                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ......................................................                                                                                                    ......................................................................                                                            ............................................................................................................................................................................                                                                                                                          ..................................................                            ................................................................................................ ......... ......... ......... ......... ......... ......... ............. ........ ........ ..... .....................................                                                                                                                                                                                                                                   ....................                                                                                                            ....................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       