















            







      




    




    ****************************************                            



    

       














































 




 





















 


 








 














 

 

 
 
   






  




 

 

 
 
   






  





















     








        












 








 



                																																	         																																																			                            																																																																																																																																																																																																																							  																																																																																																																																																																							  																																																							                                                  																																										                                                         																																																		            																			                                                                                                     																																																																										    									                                              																									                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            																																																						   																																																																																																																																																																																																																																	   									   											    																																																																																														                              																																																																																																																																																	         																                               								                     																																																																																																																																																																																																																																																																										  																								      						          																																																																																																																																																									        					          																																																																							  																																																																												            																																																																																																																																																																																																																																																																																																																																																																  																																																																					       																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																															          																																																																																																																																																																																																							**********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                    **********************                 **********************                                                     ****************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                                                                                                              


 

  


 


 


 

  


 


 























































































 

 












































 





																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								                        			                  																																																																																																																																																																																																																																																																																																																																																																																																																												                  																																																																																																																															                      ......................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 .............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................    .........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             .....................................................................................................................................................................................................................................................................              ............................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                            