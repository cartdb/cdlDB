







    



    














     














     































  





  











  







































































***************    ************************************************************************************************************************













    





  *****************



















****    ************    ****







    

****

  






















************      ********** 










 


 






    

   ****************************************************************************************************************************************************************************************    ****





 **** ********************************************* *********************************************************************************************************************  *******************  ****************  ****************************  ************









































    








































  





  



****    ********


  


  


       

   

   

   

       



    





  





  





  





  



  



  





  







***************************************************************************************************************************************************************************************************************************************************

  



    





 







     

 


 







     

 


 







    

 


 







 



 


 


 

**************************************************************************************************************************************************************                        






























*****************************************************************************************************************************************************************************************



																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				       																																																																																																																																																																																																																									            					                                																																																																																																																																																																																																																																																																																							                                																																					        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			   																																																																																																																																																			                       										         																																				 																																																																																																																																																																																																											    																																																																																																																																																																																																																																																																			                        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			     																																																																																																																																																																																																											  																																																																																																																																																																											 																																																																																																																																																																																																																																																										                                                                       																																																																																																																																																											       																																																																																																																																																																																																																																																																																																						   																																																																																																																																													   										   																																																																																																																																																																																																																																																																																																																																																																     																											    																																																																																																																																																	 																																																																																																																																																																																																																																																																																																																						 																																																																																																																																																																																																																																  															  																																																															     																																																																																																																												      																																																																																																																																																																																																											                                                         				 													   									                                                                                                     																																																												                                                                                                                                                    ..........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                  ..............................................................................................................................................................................................................................................................................................................................    ..............    ...................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   