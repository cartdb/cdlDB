    



  







    



    
                                                







                                                                    





                                                                                                                                                                                    

        














                                                                                          






                                                                                                                                                                                                                                                              



            ********

      



                        

      *****************     **                                                                















****************************************                        ****

                *****         *****                                          






























***                  

      

      

      *********************************************                                                                               *********************************************                                                                                                                   *********************************************                                                                                                                      

                     






















         






















         																																																																																																																																																																																													      																																																																																																																																																																																	 										  																																						       																																																																																																																																																																						   																																				            									                                																																																						          																																																																																																																																																																																																																											                                																																																																																																																																																																																	    																		                                																					                                           																																											                                                                                                                                                                       																														  					                          																																																								   																																																		                                                                                                       																		   								   																																																																																				                         						                                                                           						   					                																																																																																																			    																								        																				                  							                       																																																																		                        																				         													  			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             																									                                 																																																																																																																																					            																																																									    																																																																																				               							                                                                                                                                                                                     																		                          																																																																																			              						         																															                                                                																																																																						                                                             																																	         																									    																																																																																																											     																					     																											         					        																							   																																																																																								       																																																																																																																																																													       						       																						 																																					  																																																																		   																									   																																										                                			    																																																				      																																																                                           																																																																																																																																																																																																																																																																																										  																			   																							  																																																																																																																																																																																																																																																		  																																				  															      																																																																																																					      																																																																																																																																			          											                                                                                  																																																																																																																																																																																																			          									      																																																																																																																																			  																																																																																															             																																																																																																																																																																																																																																																																																							 																												                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ........................................................................................                                                                                                                                                                                                                                                                                                                                                                  ................................                                                                                                                                    .                              .                               ..                                                                                      ...................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            