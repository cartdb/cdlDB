																																																																																																																																																																																																																																	                																																																											  									               					            			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      																																						                                                                     					   																																																				                         													                                                                    																																																																																																																																																																																																										**************  ********																																																									       																	    																					****************																																																																																																																																												    														   																																																																																													                     																																																																																																																																																																																																											                                            																																																																																																																																																																																							                                  																																																																																																																																																																																																																																											           																																							      																																																		       																																																																																															    																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																						          							 																																																																																 																																																																																																																																																									 																																																																																																																																																																																																																																																																																													           									    																																							                                                                                 																																																																																																												    																																																																																																																																																																																																																																																																																																																								 				 																																	 																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			       																																																																																																																																																																																																																																																																	       																																																		                																																																																																																															             																																				      								                                																														      																																																																																																												            																																																																																																                  																																																																													


										                    																																																											                                   																																																																																																	                 																	    																																																																																									     																																																																																																																																															    																																																      																																																																																																																		                                																																																																										   																							  																																																																																																																												     																																																																																		
     																																																																																																																																																																																																																																																																																																																																																																									                   																																  																			      																																																										    																																																					        																		                                                   ................                ................                                                                                           ................                                 ......                              .........         ........................                                                                      ......                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ....................................................................................................................................................................                            .....................................................................................................................................................................................................................................................................................................................................................................................................................................................................                ....  .................................................................................................................................................                                      .............   ... ......         ... ........              ......................................                                                                                   .......  ................................................................                                               ...............................................................................................................................    ..............  ..              ..  .....................             ..............                  ............                                                        ..........                   .....................        ......................................................................                   ..............................................                                                                                                                                      ...................................................                                                                                                                                                                                                                                     ...................                             .....................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  